module fifo #(
    parameter DEPTH = 16,
    parameter WIDTH = 32
) (
    input logic clk,
    input logic rst,
    input logic [WIDTH-1:0] d_in,
    output logic [WIDTH-1:0] d_out
);

// internal logic

endmodule
