// generated
module gen_v376();
    integer j;
    initial begin
        for (j=0;j<10;j=j+1) begin
            if (j%2==0) ;
        end
    end
endmodule
