module top_mod (
    input logic a
);

module inner_mod (
    input logic b
);

endmodule

endmodule
